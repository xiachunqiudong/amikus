module decoder(
  input  wire [31:0] inst,
  output wire        instInfo,
  output wire [4:0]  lsrc1,
  output wire [4:0]  lsrc2,
  output wire [4:0]  ldst
);

  


endmodule