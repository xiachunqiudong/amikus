`define XLEN 64