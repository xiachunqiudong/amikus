module alu(
  input  wire [`XLEN-1:0] src1,
  input  wire [`XLEN-1:0] src2,
  input  wire             isAdd,
  input  wire             isSub,
  input  wire             isAnd,
  output wire [`XLEN-1:0] result
);



endmodule